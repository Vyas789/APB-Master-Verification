package apb_master_pkg;
`include "uvm_macros.svh"
 import uvm_pkg::*; 
`include"apb_master_defines.sv"
`include "apb_master_sequence_item.sv"
`include "apb_master_sequence.sv"
`include "apb_master_sequencer.sv"
`include "apb_master_driver.sv"
`include "apb_master_active_monitor.sv"
`include "apb_master_passive_monitor.sv"
`include "apb_master_active_agent.sv"
`include "apb_master_passive_agent.sv"
`include "apb_master_scoreboard.sv"
`include "apb_master_subscriber.sv"
`include "apb_master_environment.sv"
`include "apb_master_test.sv"
endpackage
